module multiplier(
    input wire mult, clk, reset,
    input wire [31:0] A,B,
    output wire[31:0] min,max
);


    
endmodule