module multiplier(
    input wire clk
    input wire reset,
    input wire mult_on,
    input wire [31:0] A,
    input wire [31:0] B,
    output wire[31:0] min
    output wire[31:0] max
);


    
endmodule