module divider(
    input wire Div,  
    input wire clk, 
    input wire reset,
    input wire SrcA, 
    input wire SrcB,
    output wire Dzero,
    output wire [31:0]min, max 
);


    
endmodule