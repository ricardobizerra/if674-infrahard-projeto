module divider(
    input wire clk, 
    input wire reset,
    input wire div_on,  
    input wire SrcA, 
    input wire SrcB,
    output wire Dzero,
    output wire [31:0]min, 
    output wire [31:0]max 
);


    
endmodule