module divider(
    input wire Div, clk, reset,
    input wire SrcA, SrcB,
    output wire Dzero,
    output wire [31:0]min, max 
);


    
endmodule